typedef uvm_sequencer # (my_transaction) my_sequencer